module half_adder(a,b,sum,carry)
sum = a^b;
carry = ab;
endmodule